module uart_tx_op_tb (
  
);

uart_rx_op .uart_rx_op_1(
  
);
endmodule //uart_tx_op_tb