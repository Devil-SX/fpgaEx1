module uart_tx_op_tb();
	clk_divider clk1(/*AutoInst*/);	
	clk_divider clk2(/*AutoInst*/);	

endmodule
